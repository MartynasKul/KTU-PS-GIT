
--KTU 2015
--Informatikos fakultetas
--Kompiuteriu katedra
--Kompiuteriu Architektura [P175B125] 
--Kazimieras Bagdonas

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is 
	port (
		RST_ROM 	: in std_logic;
		clk 		: in std_logic;
		ROM_CMD 	: in std_logic_vector(7 downto 0);	  
		ROM_Dout 	: out std_logic_vector(1 to 80)
		);
end ROM ;

architecture rtl of ROM is
	
	type memory is array (0 to 255) of std_logic_vector(1 to 80) ; 	
	
	constant ROM_CMDln : memory := (	  
--                     1         2         3         4         5         6         7         8 Dvi komentaro eilutes duoda bitu numerius   
--            12345678901234567890123456789012345678901234567890123456789012345678901234567890    (nuo 1 iki 80)
0=> "00000000000000100000000000000000000000000000000000000000000000000000000000000001",  --Ivedamas N1
1=> "00000000000000000000010000001000000000000000000000000000000000000000000000000010",  --Ivedamas N2
2=> "00000000000000000000001000000100000100000000000000000000000000000000000000000011",  --Ivedamas N3
3=> "00000000000000000000000100000010000000000000000000000000000000000000000000000100",  --Komentaro vieta
4=> "00010000000000000000000000000000000000000000000000000000000000000000000000000101",  --Komentaro vieta
5=> "00000000000000000000000000000000000000000000000000000000000000000000100000000111",  --Komentaro vieta
6=> "00000001000000000000000000000000000000000000000000010000000000000000000000001011",  --Komentaro vieta
7=> "00000000000000000000000000000000000000000000000000000000000000000001000000001001",  --Komentaro vieta
8=> "00000001000000000000000000000000000000000000000001000000000000000000000000000111",  --Komentaro vieta
9=> "00000000000000000000001000000010000000000000000000000000000000000000000000001010",  --Komentaro vieta
10=> "00000000000000000000000000000000000000000000000000000000000000000000110100000101",  --Komentaro vieta
11=> "00100001000000000000000000000000000000000000000000000010000000000000000000001100",  --Komentaro vieta
12=> "00000001000000000000000000000000000000000000000001000000000000000000000000001101",  --Komentaro vieta
13=> "01000000000000000000000000000000000000000000000000000000000000000000000000001110",  --Komentaro vieta
14=> "00000000000000000000000000000000000000000000000000000000000000000000000100001111",  --Komentaro vieta
15=> "00000000000000000000000000000000000000000000000000000000000000000010000000001111",  --Komentaro vieta
16=> "00000001000000000000000000000000000000000000000000000001000000000000000000010001",  --Komentaro vieta
17=> "00000001000000000000000000000000000000000000000000010000000000000000000000010010",  --Komentaro vieta
18=> "00000000100000000000000000000000000000000000000000000000000000000000000000010011",  --Komentaro vieta
19=> "00000001000000000000000000000000000000000000000000000010000000000000000000010100",  --Komentaro vieta
20=> "00000000000001000000000000000000000000000000000000000000000000000000000000001111",  --Komentaro vieta



	others => (others => '0') );   
	
	
	
	
begin
	process (RST_ROM, clk) 
		
	begin
		if 	RST_ROM'event and RST_ROM = '1'	 then 
			ROM_Dout <= ROM_CMDln(0);
		elsif clk'event and clk = '0' then
			ROM_Dout <= ROM_CMDln(to_integer(unsigned(ROM_CMD))); 
		end if;
		
	end process;
	
end rtl;